`timescale 1ns / 1ps

// Write First Mode

module DataMemoryRAM #(parameter DEPTH=256,ADDRESS_WIDTH=8,DATA_WIDTH=32)
   (
    input 			clk,
    input 			en,
    input 			WE,
    input [ADDRESS_WIDTH-1:0] 	addr,
    input [DATA_WIDTH-1:0] 	writedata,
    output reg [DATA_WIDTH-1:0] RD
    );

   reg [DATA_WIDTH-1:0] 	      RAM [DEPTH-1:0];

   initial
     begin
	//$readmemb("InstructionMemoryRAM.data",RAM,0,DEPTH-1);
	
RD = 32'b00000000000000000000000000000000;

RAM[0] = 32'b10010100001000000110111100101111;
RAM[1] = 32'b11011001011011011000111111110000;
RAM[2] = 32'b00000000111111111100000000111111;
RAM[3] = 32'b11111111111111111111111111111110;
RAM[4] = 32'b01110000001000001111001001111011;
RAM[5] = 32'b01001001111111100110110001110110;
RAM[6] = 32'b01010001110001000000100111110010;
RAM[7] = 32'b11111100000001001000001000100110;
RAM[8] = 32'b00100000011001110110000010011111;
RAM[9] = 32'b01101001110111010110100001010100;
RAM[10] = 32'b00010111010100001010011001110111;
RAM[11] = 32'b10011101001001111001111000100011;
RAM[12] = 32'b00111110000011011001101100100101;
RAM[13] = 32'b11000100111101001010001100101110;
RAM[14] = 32'b00111111000110100001010001011001;
RAM[15] = 32'b01010001000001011101001011001001;
RAM[16] = 32'b10110101001011100111101101111110;
RAM[17] = 32'b00001011100001101010111101000100;
RAM[18] = 32'b10111000100101110111010000000111;
RAM[19] = 32'b10000101110100001011111100101010;
RAM[20] = 32'b00111100010110100111000000010001;
RAM[21] = 32'b01010011110001000101001000010000;
RAM[22] = 32'b10110000000001000010111111011010;
RAM[23] = 32'b00110010010001111010100010101001;
RAM[24] = 32'b00010110101110000010010010000101;
RAM[25] = 32'b10010111100001111011111010101110;
RAM[26] = 32'b11110000110101011100101000011110;
RAM[27] = 32'b00010011111111001110100101010111;
RAM[28] = 32'b11010111001111000101110100001110;
RAM[29] = 32'b11010101110010111110011001111000;
RAM[30] = 32'b00101110100001101001000011101101;
RAM[31] = 32'b11001100110001010010010001011110;
RAM[32] = 32'b01110110010110010111011001010101;
RAM[33] = 32'b01000001100000110000111001110100;
RAM[34] = 32'b00010100100000100110000011111111;
RAM[35] = 32'b01000000010111110010010110001111;
RAM[36] = 32'b10010011110001000100110010000101;
RAM[37] = 32'b10000010110000000111011111110100;
RAM[38] = 32'b11001100000011110000111000000001;
RAM[39] = 32'b10101111010101001000110100101010;
RAM[40] = 32'b01100010111001011110001001011001;
RAM[41] = 32'b11111100010111000010001011001000;
RAM[42] = 32'b11000001110000100000011011001010;
RAM[43] = 32'b01001010111100100010100011101001;
RAM[44] = 32'b10000100111111111000001110110101;
RAM[45] = 32'b10100101110001010000010011111100;
RAM[46] = 32'b01000011010000000010110001111101;
RAM[47] = 32'b00101001101101001100010001010000;
RAM[48] = 32'b01111100100110111111001111001100;
RAM[49] = 32'b01100001000101011001000111110010;
RAM[50] = 32'b10000110100010100000000111011101;
RAM[51] = 32'b00101011011010000000100000010000;
RAM[52] = 32'b01000110000001011010111101001101;
RAM[53] = 32'b00100010010100001100111101110111;
RAM[54] = 32'b10111001000010000101010101010101;
RAM[55] = 32'b01110100110011010000101010111111;
RAM[56] = 32'b00001100011101100101001100111010;
RAM[57] = 32'b01010110000001000010010011011111;
RAM[58] = 32'b01010110010000011111010000111001;
RAM[59] = 32'b10000000110010101000000001011000;
RAM[60] = 32'b11011110010111000000000010101110;
RAM[61] = 32'b01110000100000000100100111100001;
RAM[62] = 32'b01001010110110111111110001000010;
RAM[63] = 32'b10000101000111000110010011111011;
RAM[64] = 32'b01111001011101011111110001101010;
RAM[65] = 32'b10100101010100010111011100110011;
RAM[66] = 32'b00010000101111110001110111011001;
RAM[67] = 32'b00000011101000100111010100010011;
RAM[68] = 32'b11110011101100101111010110000111;
RAM[69] = 32'b10111000011010001110011111111010;
RAM[70] = 32'b10100100010110111011100010100001;
RAM[71] = 32'b01100100001000110001011111011010;
RAM[72] = 32'b00000110100011111011101011111011;
RAM[73] = 32'b11010110100011011100110100000111;
RAM[74] = 32'b01010010010100001101010110111011;
RAM[75] = 32'b01001101011111110101000101111001;
RAM[76] = 32'b11010001110111010001000011111101;
RAM[77] = 32'b00011000001111011101111100000010;
RAM[78] = 32'b11101101100011010001100000001110;
RAM[79] = 32'b00010011010000100100100010001101;
RAM[80] = 32'b00000111111110001001001101111101;
RAM[81] = 32'b10100011000100110101110110001011;
RAM[82] = 32'b10110000000011111000110010001110;
RAM[83] = 32'b10100100100000010011110000110011;
RAM[84] = 32'b10111000001001101101001000101000;
RAM[85] = 32'b01111100010000111101100101010010;
RAM[86] = 32'b11010010111110001100101111111001;
RAM[87] = 32'b10000101010010001000000011111101;
RAM[88] = 32'b10111101101010100111111100010001;
RAM[89] = 32'b01111100000101101010101111111101;
RAM[90] = 32'b11001101100101110111111000101010;
RAM[91] = 32'b10001010111110011101011111111010;
RAM[92] = 32'b00110011000110000010011100011011;
RAM[93] = 32'b00101001100010010010110110000100;
RAM[94] = 32'b01111100100001101110011111000000;
RAM[95] = 32'b11100110110100011111000110100001;
RAM[96] = 32'b10001101000100011001011010000010;
RAM[97] = 32'b01000011010100010111001101111110;
RAM[98] = 32'b01011101000001010100111101010110;
RAM[99] = 32'b01110111111001100101001011111111;
RAM[100] = 32'b01110000110011010110100011100001;
RAM[101] = 32'b11001000100011010111111000110100;
RAM[102] = 32'b00010011000110011100010011110110;
RAM[103] = 32'b11111111110010101101000101001010;
RAM[104] = 32'b10011100010111110100101100010111;
RAM[105] = 32'b11010110001110001101100100001011;
RAM[106] = 32'b10001101100101100111111101111101;
RAM[107] = 32'b10100111110001001100010001000011;
RAM[108] = 32'b10111001011001110100001011001110;
RAM[109] = 32'b11111001110101100100110001000000;
RAM[110] = 32'b10100101000011010011010000010111;
RAM[111] = 32'b10011001001101001101000100011100;
RAM[112] = 32'b10100110001011000001000100001000;
RAM[113] = 32'b10011101111010010001000100110111;
RAM[114] = 32'b11110101001100100111010011000110;
RAM[115] = 32'b10111110101100010100100010010011;
RAM[116] = 32'b00000101011001100101100010010101;
RAM[117] = 32'b00100110000010001011111001101111;
RAM[118] = 32'b10111010100001011000100111000110;
RAM[119] = 32'b00111110100111001110110010111011;
RAM[120] = 32'b11100001000110001110011110100001;
RAM[121] = 32'b11111100001111000111000101100101;
RAM[122] = 32'b01101101010110111001010000101100;
RAM[123] = 32'b01010000111011011000110011000001;
RAM[124] = 32'b10000100000110001100010101111001;
RAM[125] = 32'b00111111111001110110001111001011;
RAM[126] = 32'b00000111100101000111100010100000;
RAM[127] = 32'b10101010101010101010101010101010;
RAM[128] = 32'b10110100001100110000100001111110;
RAM[129] = 32'b10110110101101101111111001100101;
RAM[130] = 32'b10011111010001111000100010011000;
RAM[131] = 32'b00001111010011001000010110001001;
RAM[132] = 32'b00100010011101111100001110100011;
RAM[133] = 32'b01101011000011001001001100100111;
RAM[134] = 32'b00111011011111001010001011110000;
RAM[135] = 32'b10100011000100111011110001101000;
RAM[136] = 32'b01000110001000110111011001011001;
RAM[137] = 32'b10110110100101110000100110000010;
RAM[138] = 32'b10111110110001111110101001010111;
RAM[139] = 32'b00011101001010101101111100001111;
RAM[140] = 32'b01110100111010011000110110010100;
RAM[141] = 32'b11110001111111011010110100001000;
RAM[142] = 32'b01001001110010100111010010001011;
RAM[143] = 32'b01111100100000001101000110001111;
RAM[144] = 32'b00010111111011001001101001010100;
RAM[145] = 32'b11110001111110100111101011110010;
RAM[146] = 32'b10110000101000000001011011111110;
RAM[147] = 32'b11101100111111011010100011000100;
RAM[148] = 32'b01011000110000000101100110101000;
RAM[149] = 32'b10100111011111110100101000000000;
RAM[150] = 32'b01001111010101010111100000011011;
RAM[151] = 32'b11001101001101000100100100010111;
RAM[152] = 32'b11000011000000101100101100101000;
RAM[153] = 32'b10010000001000111110011010100111;
RAM[154] = 32'b11111110000001011111011110001110;
RAM[155] = 32'b00100100100000110100010100111101;
RAM[156] = 32'b11110110000001100110010011000010;
RAM[157] = 32'b11100100100111000101001101101001;
RAM[158] = 32'b10101100111001010100111110001010;
RAM[159] = 32'b00011110011001110110111011000010;
RAM[160] = 32'b01000100011110010111011001001110;
RAM[161] = 32'b11010001010110011000110110000101;
RAM[162] = 32'b00001011110110010111011111010000;
RAM[163] = 32'b11001011110110001110001111110111;
RAM[164] = 32'b00100011110010011011001000101110;
RAM[165] = 32'b10010101011110010100010010011110;
RAM[166] = 32'b11110100011010111101101001110011;
RAM[167] = 32'b10010010010111101100110010110110;
RAM[168] = 32'b11110100001100111111111010101001;
RAM[169] = 32'b01000000111101010101011001011001;
RAM[170] = 32'b11101100101111010111001011011000;
RAM[171] = 32'b10011110111000111001110000110010;
RAM[172] = 32'b00111000110011100101001001101001;
RAM[173] = 32'b01010011011110011001011000011101;
RAM[174] = 32'b01101001011101011011101011100011;
RAM[175] = 32'b10101101110100010101011101111000;
RAM[176] = 32'b11001010111111011001100011101100;
RAM[177] = 32'b00011110000100011100100011000011;
RAM[178] = 32'b01011001001001110101101001101010;
RAM[179] = 32'b10100100111000110101000011011010;
RAM[180] = 32'b00100101011001100010010101011101;
RAM[181] = 32'b01100110110100100010011000011001;
RAM[182] = 32'b11111110011010010110111111101100;
RAM[183] = 32'b11100000110111010001111000011010;
RAM[184] = 32'b00000011110001011000110110011111;
RAM[185] = 32'b10110000010000110011110110001110;
RAM[186] = 32'b11101001100111011111010100011101;
RAM[187] = 32'b01101110111011000110010010011000;
RAM[188] = 32'b11010111110000011011110110010011;
RAM[189] = 32'b11010001101100010011110110010101;
RAM[190] = 32'b01001100111010110011110000101001;
RAM[191] = 32'b10001001111110011110111100110111;
RAM[192] = 32'b01111100111000011110001011010110;
RAM[193] = 32'b00010011011011100011101011100000;
RAM[194] = 32'b10111101011110110001101011001100;
RAM[195] = 32'b10101111100001110001001110101010;
RAM[196] = 32'b00110001101110010100100001011111;
RAM[197] = 32'b00001010001000111010010010100000;
RAM[198] = 32'b10001101111111001001101010110111;
RAM[199] = 32'b11100101110001111100011110001110;
RAM[200] = 32'b01100111010101010100011011000100;
RAM[201] = 32'b01010101100110101100000110101100;
RAM[202] = 32'b11110101001110101001000101100001;
RAM[203] = 32'b11110110000101111001001110110111;
RAM[204] = 32'b00101011010000100110101010111011;
RAM[205] = 32'b00000110000001000001001100101011;
RAM[206] = 32'b01100100101111111100111010000100;
RAM[207] = 32'b11010001010101001000110100100111;
RAM[208] = 32'b11010010110010001000111111010101;
RAM[209] = 32'b01101011111011001110000110101111;
RAM[210] = 32'b00000110000111000100101100110010;
RAM[211] = 32'b11010110101011010110101010110011;
RAM[212] = 32'b10111011011100011110000100000100;
RAM[213] = 32'b11111100011010101011010010100101;
RAM[214] = 32'b01010010011110001101000011010000;
RAM[215] = 32'b11101101011101110100000110010010;
RAM[216] = 32'b11010000011000100110011101101001;
RAM[217] = 32'b10011011001010111011101110000010;
RAM[218] = 32'b11100110100001111011000100001100;
RAM[219] = 32'b10011110111110001111101101010011;
RAM[220] = 32'b01010101110011000000011001000100;
RAM[221] = 32'b10010011111001111111000000001000;
RAM[222] = 32'b10010101010101000110110110111010;
RAM[223] = 32'b01110101000010011010110101011110;
RAM[224] = 32'b10111101001100110001000010110011;
RAM[225] = 32'b00011101111010110110110101001111;
RAM[226] = 32'b11000000010111111000101101110011;
RAM[227] = 32'b01000000101000110110011001111001;
RAM[228] = 32'b00000001111101000100000110000000;
RAM[229] = 32'b10010011000010000100111011010001;
RAM[230] = 32'b00011101011111110001111010110101;
RAM[231] = 32'b00010000111101011000000101001011;
RAM[232] = 32'b01000001100111001101100110100111;
RAM[233] = 32'b01101000000110111100111011100010;
RAM[234] = 32'b00110100101100001000101110110010;
RAM[235] = 32'b00011011010010010110101000110010;
RAM[236] = 32'b11101111010110001000010111010111;
RAM[237] = 32'b11100100001000000000111001101010;
RAM[238] = 32'b11010010010110110111011100111110;
RAM[239] = 32'b00000101010111000011110111100010;
RAM[240] = 32'b01010101000111111100001100001111;
RAM[241] = 32'b01000010000111100100010000011101;
RAM[242] = 32'b11111100101010000000100100010101;
RAM[243] = 32'b00011010010010010011111101100110;
RAM[244] = 32'b11000100000000101100011000010111;
RAM[245] = 32'b11011011101101010010111111011010;
RAM[246] = 32'b11101000010100000011100011001100;
RAM[247] = 32'b01110100001100100011011001010100;
RAM[248] = 32'b01000010001001001110010100011010;
RAM[249] = 32'b11011101011001100001100000101000;
RAM[250] = 32'b00010010100001000011011000011011;
RAM[251] = 32'b11011111011011011001101100010001;
RAM[252] = 32'b11010100110001111100110010100010;
RAM[253] = 32'b10111100000011101110010010000101;
RAM[254] = 32'b11010010100011100010110010010001;
RAM[255] = 32'b11011010011100000111011000100010;
     end // initial begin
   
   always @(posedge clk)
     begin
	if(en)	    
	  begin
	     if(WE)
	       begin
		  RAM[addr]<=writedata;
		  RD<=writedata;
	       end
	     else
	       RD<=RAM[addr];
	     
	  end // if (en)
     end // always @ (posedge clk)
   
endmodule // DataMemoryRAM
