`timescale 1ns / 1ps

// Read First Mode

module InstructionMemoryRAM #(parameter DEPTH=256,ADDRESS_WIDTH=8,WIDTH=32)
   (
    input 			clk,
    input 			en_,
    input 			CLR,
    input [ADDRESS_WIDTH-1:0] 	addr,
    output reg [WIDTH-1:0] InstrD
    );

   reg [WIDTH-1:0] 	      RAM [DEPTH-1:0];
	
	parameter R     = 6'h00;
//	parameter NULL  = 5'h00;
	
	parameter ADD   = 6'h20;
   parameter AND   = 6'h24;
   parameter OR    = 6'h25;
   parameter SEQ   = 6'h28;
   parameter SLE   = 6'h2c;
   parameter SLL   = 6'h04;
   parameter SLT   = 6'h2a;
   parameter SNE   = 6'h29;
   parameter SRA   = 6'h07;
   parameter SRL   = 6'h06;
   parameter SUB   = 6'h22;
   parameter XOR   = 6'h26;
   
   parameter J     = 6'h02;
   parameter JAL   = 6'h03;
   
   parameter ADDI  = 6'h08;
   parameter ANDI  = 6'h0c;
   parameter BEQZ  = 6'h04;
   parameter BNEZ  = 6'h05;
   parameter JALR  = 6'h13;
   parameter JR    = 6'h12;
   parameter LHI   = 6'h0f;
   parameter LW    = 6'h23;
   parameter ORI   = 6'h0d;
   parameter SEQI  = 6'h18;
   parameter SLEI  = 6'h1c;
   parameter SLLI  = 6'h14;
   parameter SLTI  = 6'h1a;
   parameter SNEI  = 6'h19;
   parameter SRAI  = 6'h17;
   parameter SRLI  = 6'h16;
   parameter SUBI  = 6'h0a;
   parameter SW    = 6'h2b;
   parameter XORI  = 6'h0e;
   
	initial
     begin
	$readmemb("/home/sumit/ISEProjects/MIPS_CPU/src/InstructionMemoryRAM.txt",RAM);
InstrD = 32'b00000000000000000000000000000000;

//RAM[0]  ={ORI  ,5'd0 ,5'd1 ,16'b0000000000001010};
//RAM[1]  ={SW   ,5'd1 ,5'd1 ,16'b0000000000000000};
//RAM[2]  ={R    ,5'd2 ,5'd1 ,5'd2 ,5'd00,  ADD};
//RAM[3]  ={SUBI ,5'd1 ,5'd1 ,16'b0000000000000001};
//RAM[4]  ={BNEZ ,5'd1 ,5'd0 ,16'b1111111111111100};
//RAM[5]  ={6'h00,5'd00,5'd00,5'd00,5'd00,6'h00};
//RAM[6]  ={6'h00,5'd00,5'd00,5'd00,5'd00,6'h00};
//RAM[7]  ={6'h00,5'd00,5'd00,5'd00,5'd00,6'h00};
//RAM[8]  ={6'h00,5'd00,5'd00,5'd00,5'd00,6'h00};
//RAM[9]  ={6'h00,5'd00,5'd00,5'd00,5'd00,6'h00};
//RAM[10] ={6'h00,5'd00,5'd00,5'd00,5'd00,6'h00};
//RAM[11] ={6'h00,5'd00,5'd00,5'd00,5'd00,6'h00};
//RAM[12] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[13] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[14] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[15] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[16] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[17] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[18] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[19] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[20] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[21] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[22] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[23] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[24] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[25] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[26] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[27] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[28] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[29] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[30] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[31] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[32] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[33] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[34] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[35] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[36] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[37] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[38] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[39] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[40] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[41] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[42] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[43] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[44] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[45] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[46] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[47] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[48] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[49] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[50] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[51] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[52] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[53] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[54] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[55] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[56] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[57] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[58] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[59] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[60] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[61] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[62] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[63] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[64] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[65] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[66] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[67] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[68] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[69] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[70] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[71] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[72] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[73] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[74] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[75] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[76] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[77] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[78] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[79] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[80] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[81] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[82] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[83] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[84] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[85] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[86] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[87] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[88] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[89] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[90] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[91] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[92] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[93] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[94] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[95] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[96] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[97] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[98] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[99] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[100] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[101] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[102] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[103] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[104] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[105] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[106] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[107] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[108] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[109] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[110] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[111] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[112] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[113] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[114] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[115] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[116] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[117] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[118] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[119] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[120] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[121] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[122] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[123] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[124] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[125] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[126] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[127] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[128] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[129] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[130] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[131] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[132] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[133] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[134] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[135] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[136] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[137] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[138] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[139] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[140] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[141] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[142] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[143] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[144] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[145] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[146] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[147] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[148] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[149] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[150] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[151] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[152] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[153] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[154] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[155] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[156] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[157] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[158] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[159] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[160] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[161] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[162] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[163] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[164] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[165] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[166] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[167] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[168] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[169] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[170] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[171] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[172] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[173] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[174] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[175] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[176] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[177] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[178] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[179] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[180] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[181] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[182] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[183] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[184] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[185] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[186] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[187] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[188] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[189] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[190] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[191] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[192] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[193] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[194] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[195] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[196] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[197] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[198] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[199] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[200] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[201] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[202] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[203] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[204] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[205] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[206] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[207] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[208] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[209] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[210] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[211] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[212] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[213] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[214] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[215] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[216] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[217] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[218] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[219] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[220] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[221] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[222] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[223] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[224] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[225] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[226] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[227] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[228] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[229] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[230] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[231] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[232] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[233] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[234] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[235] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[236] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[237] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[238] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[239] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[240] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[241] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[242] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[243] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[244] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[245] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[246] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[247] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[248] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[249] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[250] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[251] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[252] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[253] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[254] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
//RAM[255] ={6'h00,5'h00,5'h00,5'h00,5'h00,6'h00};
     end
   
   always @(posedge clk)
		begin
			if(~en_)	    
			  begin
			     if(CLR)
                               InstrD<=0;
			     else
                               InstrD<=RAM[addr];
			  end
		end
   
endmodule // InstructionMemoryRAM
