`timescale 1ns / 1ps

// Read First Mode

module RegisterFile #(parameter NO_OF_REG=32,REG_ADDRESS_WIDTH=5,WIDTH=32)
   (
    input 			  clk,
    input 			  WE3,
    input [REG_ADDRESS_WIDTH-1:0] A1,
    input [REG_ADDRESS_WIDTH-1:0] A2,
    input [REG_ADDRESS_WIDTH-1:0] A3,
    input [WIDTH-1:0] 	  WD3,
    output [WIDTH-1:0] 	  RD1,
    output [WIDTH-1:0] 	  RD2
    );

   reg [WIDTH-1:0] 	      REG [NO_OF_REG-1:0];
   

   initial
     begin
	REG[0] = 32'b00000000000000000000000000000000;
	REG[1] = 32'b00000000000000000000000000000000;
	REG[2] = 32'b00000000000000000000000000000000;
	REG[3] = 32'b00000000000000000000000000000000;
	REG[4] = 32'b00000000000000000000000000000000;
	REG[5] = 32'b00000000000000000000000000000000;
	REG[6] = 32'b00000000000000000000000000000000;
	REG[7] = 32'b00000000000000000000000000000000;
	REG[8] = 32'b00000000000000000000000000000000;
	REG[9] = 32'b00000000000000000000000000000000;
	REG[10] = 32'b00000000000000000000000000000000;
	REG[11] = 32'b00000000000000000000000000000000;
	REG[12] = 32'b00000000000000000000000000000000;
	REG[13] = 32'b00000000000000000000000000000000;
	REG[14] = 32'b00000000000000000000000000000000;
	REG[15] = 32'b00000000000000000000000000000000;
	REG[16] = 32'b00000000000000000000000000000000;
	REG[17] = 32'b00000000000000000000000000000000;
	REG[18] = 32'b00000000000000000000000000000000;
	REG[19] = 32'b00000000000000000000000000000000;
	REG[20] = 32'b00000000000000000000000000000000;
	REG[21] = 32'b00000000000000000000000000000000;
	REG[22] = 32'b00000000000000000000000000000000;
	REG[23] = 32'b00000000000000000000000000000000;
	REG[24] = 32'b00000000000000000000000000000000;
	REG[25] = 32'b00000000000000000000000000000000;
	REG[26] = 32'b00000000000000000000000000000000;
	REG[27] = 32'b00000000000000000000000000000000;
	REG[28] = 32'b00000000000000000000000000000000;
	REG[29] = 32'b00000000000000000000000000000000;
	REG[30] = 32'b00000000000000000000000000000000;
	REG[31] = 32'b00000000000000000000000000000000;
     end // initial begin
   
   always @(negedge clk)
     begin
	if(WE3)
	  REG[A3]=WD3;
	//read_A1<=A1;
	//read_A2<=A2;
     end
   
   assign   RD1=REG[A1];
   assign   RD2=REG[A2];
   
endmodule // RegisterFile
